`timescale 1ns / 1ps

module sdramController(
  input logic clk, rst_n,
  input  logic        instr_enable,
  output logic        instr_valid,
  input  logic [24:0] instr_addr,
  output logic [31:0] instr_result,

  input  logic         data_enable,
  output logic         data_valid,
  input logic  [1:0]   data_oplen,
  input logic          data_unsigned,
  input logic  [24:0]  data_addr,
  input logic  [31:0]  data_wdata,
  input logic          data_rw,
  output logic [31:0]  data_result,

  output logic        s_clk,   output logic        s_cs_n,
  output logic        s_ras_n, output logic        s_cas_n,
  output logic        s_we_n,  output logic        s_cke,
  output logic [1:0]  s_dqm,   output logic [12:0] s_addr,
  output logic [1:0]  s_bs,    inout  logic [15:0] s_dq
);

module sextender_m(input logic [31:0]in, input logic usgn,
                 input logic [1:0]len, output logic [31:0]out);
  always_comb begin
    if (usgn) begin
      unique case (len)
        2'b00: out = { {24{1'b0}}, in[7:0] } ;
        2'b01: out = { {24{1'b0}}, in[15:0] } ;
        2'b10: out = { {24{1'b0}}, in[23:0] } ;
        2'b11: out = { in[31:0] } ;
      endcase
    end else begin
      unique case (len)
        2'b00: out = { {24{in[7]}}, in[7:0] } ;
        2'b01: out = { {24{in[15]}}, in[15:0] } ;
        2'b10: out = { {24{in[23]}}, in[23:0] } ;
        2'b11: out = { in[31:0] } ;
      endcase
    end
  end
endmodule

logic [31:0]internal_data_result;
sextender_m sextender(
  .in(internal_data_result), .usgn(data_unsigned),
  .len(data_oplen), .out(data_result));

assign s_clk = clk;

logic [3:0]startupStep;
logic [15:0]dq;
assign s_dq = dq;

logic [15:0]instr_read_delay;
logic [15:0]data_read_delay;

logic [31:0]ops[30];
logic [31:0]shittyram[100];
always_ff @(posedge clk) begin
  if (!rst_n) begin
ops[0] <= 32'h00100093;
ops[1] <= 32'h00100113;
ops[2] <= 32'h00000513;
ops[3] <= 32'h02000593;
ops[4] <= 32'h00450513;
ops[5] <= 32'h002081b3;
ops[6] <= 32'h00010093;
ops[7] <= 32'h00018113;
ops[8] <= 32'h00152023;
ops[9] <= 32'hfeb516e3;

    instr_valid <= 1'b0;
    instr_read_delay <= 16'h00;
    data_valid <= 1'b0;
    data_read_delay <= 16'h00;
  end else begin
    // TODO: Handle non aligned reads
    data_valid <= 1'b0;
    instr_valid <= 1'b0;
    if (data_enable && !data_valid && data_read_delay == 16'h00) begin
      if (data_rw) begin
        unique case (data_oplen)
          2'b00: shittyram[data_addr >> 2][7:0] <= data_wdata[7:0];
          2'b01: shittyram[data_addr >> 2][15:0] <= data_wdata[15:0];
          2'b10: shittyram[data_addr >> 2][23:0] <= data_wdata[23:0];
          2'b11: shittyram[data_addr >> 2][31:0] <= data_wdata[31:0];
        endcase
      end else begin
        unique case (data_oplen)
          2'b00:internal_data_result <= {24'h0000, shittyram[data_addr >> 2][7:0]};
          2'b01:internal_data_result <= {16'h0000, shittyram[data_addr >> 2][15:0]};
          2'b10:internal_data_result <= {8'h0000, shittyram[data_addr >> 2][23:0]};
          2'b11:internal_data_result <= {shittyram[data_addr >> 2][31:0]};
        endcase
      end
      data_read_delay <= 8;
    end else if (data_read_delay > 0) begin
      data_valid <= 1'b0;
      data_read_delay <= data_read_delay - 1;
      if (data_read_delay == 1) begin
        data_valid <= 1'b1;
        if (instr_enable) begin instr_valid <= 1'b0; end
      end
    end else if (instr_enable && !instr_valid && instr_read_delay == 16'h00) begin
      if ((instr_addr >> 2) > 18) begin $stop(); end
      instr_result <= {ops[instr_addr >> 2][31:0]};
      instr_read_delay <= 8;
      instr_valid <= 1'b0;
    end else if (instr_read_delay > 0) begin
      instr_valid <= 1'b0;
      instr_read_delay <= instr_read_delay - 1;
      if (instr_read_delay == 1) begin
        instr_valid <= 1'b1;
      end
    end
  end
end

/*
 * StartUp
 *
 * WaitStart, Precharge, Mode Register State
 * AutoRefresh 1-8,
 *
 */


/*
logic [6:0]powerupState;
localparam logic[6:0] MAX_POWERUP_STATE = 7'd80;
localparam logic[15:0] HI_Z = 16'hZZZZ;

always_ff @(posedge clk) begin
  if (!rst_n) begin
    powerupState <= 7'h00;
  end else begin
    if (powerupState <= MAX_POWERUP_STATE) begin
      powerupState <= powerupState + 1;
    end
  end
end

task automatic nop;
  begin
    s_cke   <= 1;
    s_cs_n  <= 0;
    s_ras_n <= 1;
    s_cas_n <= 1;
    s_we_n  <= 1;
    s_dqm   <= 0;
    s_bs    <= 0;
    s_addr  <= 0;
    dq    <= HI_Z;
  end
endtask

task precharge_bank_0;
  input [1 : 0] dqm_in;
  input [15 : 0] dq_in;
  begin
    cke   = 1;
    cs_n  = 0;
    ras_n = 0;
    cas_n = 1;
    we_n  = 0;
    dqm   = dqm_in;
    ba    = 0;
    addr  = 0;
    dq    = dq_in;
  end
endtask

task precharge_bank_1;
  input [1 : 0] dqm_in;
  input [15 : 0] dq_in;
  begin
    cke   = 1;
    cs_n  = 0;
    ras_n = 0;
    cas_n = 1;
    we_n  = 0;
    dqm   = dqm_in;
    ba    = 1;
    addr  = 0;
    dq    = dq_in;
  end
endtask

task automatic precharge_banks;
  begin
    s_cke   <= 1;
    s_cs_n  <= 0;
    s_ras_n <= 0;
    s_cas_n <= 1;
    s_we_n  <= 0;
    s_dqm   <= 0;
    s_bs    <= 0;
    s_addr  <= 1024; // A10 = 1
    dq    <= HI_Z;
  end
endtask

task automatic auto_refresh;
  begin
    s_cke   <= 1;
    s_cs_n  <= 0;
    s_ras_n <= 0;
    s_cas_n <= 0;
    s_we_n  <= 1;
    s_dqm   <= 0;
    s_bs    <= 0;
    s_addr  <= 0;
    dq    <= HI_Z;
  end
endtask

task automatic load_mode_reg;
  input [12 : 0] op_code;
  begin
    s_cke   <= 1;
    s_cs_n  <= 0;
    s_ras_n <= 0;
    s_cas_n <= 0;
    s_we_n  <= 0;
    s_dqm   <= 0;
    s_bs    <= 0;
    s_addr  <= op_code;
    dq    <= HI_Z;
  end
endtask


task automatic bank_active;
  input [ 1 : 0] bank;
  input [12 : 0] row;
  begin
    s_cke   <= 1;
    s_cs_n  <= 0;
    s_ras_n <= 0;
    s_cas_n <= 1;
    s_we_n  <= 1;
    s_dqm   <= 0;
    s_bs    <= bank;
    s_addr  <= row;
    dq    <= HI_Z;
  end
endtask

task automatic write;
  input [ 1 : 0] bank;
  input [ 8 : 0] column;
  input [15 : 0] dq_in;
  begin
    s_cke   <= 1;
    s_cs_n  <= 0;
    s_ras_n <= 1;
    s_cas_n <= 0;
    s_we_n  <= 0;
    s_dqm   <= 0;
    s_bs    <= bank;
    s_addr  <= column;
    dq    <= dq_in;
  end
endtask

task automatic read;
  input [ 1 : 0] bank;
  input [ 8 : 0] column;
  begin
    s_cke   <= 1;
    s_cs_n  <= 0;
    s_ras_n <= 1;
    s_cas_n <= 0;
    s_we_n  <= 1;
    s_dqm   <= 0;
    s_bs    <= bank;
    s_addr  <= column;
    dq    <= HI_Z;
  end
endtask

always_ff @(posedge clk) begin
  if (!rst_n) begin
    result <= 32'h0000;
  end else begin
    case (powerupState)
      'd1: nop;  //0-8 Nop
      'd9: precharge_banks;  //9 Precharge ALL Bank
      'd10: nop;  //10-11 Nop, tRP's minimum value is 20ns
      'd12: auto_refresh;  //12 Auto Refresh
      'd13: nop;  //13-20 Nop, tRFC's minimum value is 66ns
      'd21: auto_refresh;  //21 Auto Refresh
      'd22: nop;  //22-29 Nop, tRFC's minimum value is 66ns
      'd30: load_mode_reg(13'b0001000100011);  //30 Load Mode: Lat = 2, BL = 8, Seq
      'd31: nop;  //31 Nop, 2tCLK
      'd33: bank_active(0, 0);  //33 Active: Bank = 0, Row = 0
      'd34: nop;  //34-35 Nop
      'd36: write(0, 200, result + 1);  //36 Write : Bank = 0, Col = 200
      'd37: begin result <= 32'h0000; nop; end  //37 Nop
      'd38: nop;  //38 Nop
      'd39: nop;  //39-40 Nop
      'd50: bank_active(0, 0);  //50 Active: Bank = 0, Row = 0
      'd51: nop;  //51-52 Nop
      'd53: read(0, 200);  //53 Read Bank = 0, Col = 200
      'd54: nop;  //54 Nop
      'd55: nop;
      'd56: result <= {16'h00, s_dq};  //55 Nop
      default:;
    endcase
  end
end*/

endmodule
