module fakeram(
  input logic clk, rst_n,
  input logic [31:0]addr,
  input logic [31:0]val,
  input logic rw,
  output logic [31:0]res
  );

  logic [31:0]cram[1024];

  initial begin
    integer i;
    for (i = 0; i < 1024; i += 1) begin
      cram[i] <= 32'h0000;
    end
    for (i = 0; i < 64; i += 1) begin
      cram[i] <= i;
    end
    cram[ 0] <= 32'b0000000_00000_00000_000_00000_0110011; /// NOP
    cram[ 1] <= 32'b0000000_00000_00000_000_00000_0110011; /// NOP
    cram[ 2] <= 32'b0000000_00000_00000_000_00000_0110011; /// NOP
    cram[ 3] <= 32'b000010000001_00010_000_00010_0010011 ; /// x2 = x2 + 0x41
    cram[ 4] <= 32'b000000100001_00000_000_00001_0010011 ; /// x1 = x0 + 0x21
    cram[ 5] <= 32'b1111111_00001_00010_010_11111_0100011; /// sw x1, (-1)x2
    cram[ 6] <= 32'b111111111111_00010_010_00011_0000011 ; /// lw x3, (-1)x2
    cram[ 7] <= 32'b01010101010101010101_00100_0110111   ; /// x4 = 0x0101 << 12
    cram[ 8] <= 32'b010101010101_00100_000_00100_0010011 ; /// x4 = x0 + 0x01
    cram[ 9] <= 32'b01010101010101010101_00100_0010111   ; /// x4 = 0x0101 << 12 + pc
    cram[10] <= 32'b0000000_00011_00001_100_00001_0110011; /// x1 = x1 ^ x3
    cram[11] <= 32'b0000000_00011_00001_100_00011_0110011; /// x3 = x2 ^ x3
    cram[12] <= 32'b0000000_00011_00001_100_00001_0110011; /// x1 = x1 ^ x3
    cram[13] <= 32'b000000000000_00000_000_00001_0010011 ; /// x1 = 0
    cram[14] <= 32'b000000010000_00000_000_00010_0010011 ; /// x2 = 16
    cram[15] <= 32'b000000000001_00001_000_00001_0010011 ; /// x1 = x1 + 1
    cram[16] <= 32'b1111111_00010_00001_001_11001_1100011; /// bne x1, x2, -8
    cram[17] <= 32'b111111111111_00000_000_00001_0010011 ; /// x1 = 0
    cram[18] <= 32'b0000000_00000_00000_000_00000_0110011; /// NOP
    cram[19] <= 32'b0000000_00000_00000_000_00000_0110011; /// NOP
    cram[20] <= 32'b0000000_00000_00000_000_00000_0110011; /// NOP
  end

  always @(clk) begin
    if (clk) begin
      if (addr == 32'h60) begin $stop; end
      if (rw) begin
        res <= cram[addr >> 2];
      end
    end else begin
      if (!rw) begin
        cram[addr >> 2] <= val;
      end
    end
  end
endmodule
